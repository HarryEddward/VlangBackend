module main

import fmt

// Función principal
fn main() {
    mut edad := 25
	var nombre string = "adrian"

	println("$nombre: $edad")
}
